<HTML><HEAD><TITLE>OpenGL - Demos</TITLE></HEAD><BODY><CENTER>

<A HREF="../progs.html"><IMG SRC="../opengl.jpg"></A><BR>

<H1><A HREF="./">demos/</H1></A>

<BR><IMG SRC="../divider.gif"><BR>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="atlantis.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Swimming around with sharks, dolphins and whales.<BR>
  <BR> Source code: <A HREF="atlantis/">source directory</A>.<BR>
  <BR> Executable: <A HREF="atlantis/atlantis.exe">atlantis.exe</A>.<BR>
  <BR> Snapshots: <A HREF="atlantis.jpg">fish (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="chess.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Classical chess game with a crazy twist.<BR>
  <BR> Source code: <A HREF="chess/">source directory</A>.<BR>
  <BR> Executable: <A HREF="chess.bat">chess.bat</A>.<BR>
  <BR> Snapshots: <A HREF="chess.jpg">in game (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="geoface.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Contort this face as much as you want.<BR>
  <BR> Source code: <A HREF="geoface/">source directory</A>.<BR>
  <BR> Executable: <A HREF="geoface.bat">geoface.bat</A>.<BR>
  <BR> Snapshots: <A HREF="geoface.jpg">smile (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="glutmech.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Walking (but not talking) vulcan gunner.<BR>
  <BR> Source code: <A HREF="glutmech/glutmech.c">glutmech.c</A>.<BR>
  <BR> Executable: <A HREF="glutmech/glutmech.exe">glutmech.exe</A>.<BR>
  <BR> Snapshots: <A HREF="glutmech.jpg">shaded (shown)</A>, <A HREF="glutmech1.jpg">walking</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="ideas.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> The classic SGI demonstration program.<BR>
  <BR> Source code: <A HREF="ideas/">source directory</A>.<BR>
  <BR> Executable: <A HREF="ideas/ideas.exe">ideas.exe</A>.<BR>
  <BR> Snapshots: <A HREF="ideas.jpg">shadow (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="opengl_logo.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Cool OpenGL logo that spins into place.<BR>
  <BR> Source code: <A HREF="opengl_logo/">source directory</A>.<BR>
  <BR> Executable: <A HREF="opengl_logo/opengl_logo.exe">opengl_logo.exe</A>.<BR>
  <BR> Snapshots: <A HREF="opengl_logo.jpg">final (shown)</A>, <A HREF="opengl_logo1.jpg">motion</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="rollercoaster.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Excellent rollercoaster simulation (you can really feel this one!).<BR>
  <BR> Source code: <A HREF="rollercoaster/">source directory</A>.<BR>
  <BR> Executable: <A HREF="rollercoaster.bat">rollercoaster.bat</A>.<BR>
  <BR> Snapshots: <A HREF="rollercoaster.jpg">cart (shown)</A>, <A HREF="rollercoaster1.jpg">rush</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="underwater.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Caustic effects as viewed in underwater scenes.<BR>
  <BR> Source code: <A HREF="underwater/">source directory</A>.<BR>
  <BR> Executable: <A HREF="underwater.bat">underwater.bat</A>.<BR>
  <BR> Snapshots: <A HREF="underwater.jpg">greenish sea (shown)</A>, <A HREF="underwater1.jpg">cube underwater</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="walker.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Walking motion simulator (customizable).<BR>
  <BR> Source code: <A HREF="walker/">source directory</A>.<BR>
  <BR> Executable: <A HREF="walker/walker.exe">walker.exe</A>.<BR>
  <BR> Snapshots: <A HREF="walker.jpg">walk (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR>
<TABLE BORDER=3 WIDTH=520 CELLPADDING=6>
<TR>
 <TD><IMG SRC="yacme.jpg"></TD>
 <TD VALIGN=TOP>
  <BR> Color editor with a very nice interface.<BR>
  <BR> Source code: <A HREF="yacme/">source directory</A>.<BR>
  <BR> Executable: <A HREF="yacme/Editor.exe">yacme.exe</A>.<BR>
  <BR> Snapshots: <A HREF="yacme.jpg">default (shown)</A>.<BR>
 </TD>
</TR>
</TABLE>

<BR><IMG SRC="../divider.gif"><BR>

<H5>Copyright &copy; 1997 Silicon Graphics Incorporated.</H5>

</CENTER></BODY></HTML>
